module psdsqrt
      #(parameter NBITSIN = 32) (
        input clock,
				input reset,
				input start,
				input stop,
				input [NBITSIN-1:0] xin,
				output reg [NBITSIN/2-1:0] sqrt
			  );



endmodule
