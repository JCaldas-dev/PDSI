`timescale 1ns / 1ns

module reg_bank_tb;